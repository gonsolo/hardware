module laber;

initial begin
	$display("laber laber");
end

hurz hurz_instance();
endmodule

