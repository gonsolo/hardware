module nille(
	x
);
input x;

initial begin
	$display("nille");
end

endmodule

