module laber;

initial begin
	$display("laber laber");
end

hurz hurz1();

endmodule

