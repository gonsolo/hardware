module laber;

initial begin
	$display("laber laber");
	$finish;
end

//hurz hurz1();


endmodule

