module laber(
	clk
);
input clk;

nille nille1(clk);

initial begin
	$display("Initializing laber");
	$finish;
end

//hurz hurz1();

endmodule

