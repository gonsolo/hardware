module nille(
	clk
);
input clk;

initial begin
	$display("Initializing nille");
end

endmodule

